LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.all;
ENTITY run_modelsim IS
	PORT(
		FREQUENCY: IN STD_LOGIC_VECTOR(22 DOWNTO 0);
		CLK :IN STD_LOGIC;
		RST: IN STD_LOGIC;
		PHASE: OUT STD_LOGIC_VECTOR(22 DOWNTO 0)
	);
END run_modelsim;

ARCHITECTURE arch_run_modelsim  OF run_modelsim IS
	

BEGIN

END ARCHITECTURE;